module counter_days (
    input clk,
    input rst_n,
    input mode_day,
    input up,
    input down,
    input tick_day,
    input [5:0] max_days,
	 output ok
);

    assign ok = rst_n; 

endmodule 